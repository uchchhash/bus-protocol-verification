package i2c_m_agnt_pkg;

  //----- Include UVM Macros -----//
  `include "uvm_macros.svh"

  //----- Include Agent Package classes -----//
  `include "i2c_m_sequence_item.sv"
  `include "i2c_m_sequence_base.sv"
  `include "i2c_m_sequence_lib.sv"	

  `include "i2c_m_agent_config.sv"
  `include "i2c_m_monitor.sv"
  `include "i2c_m_driver.sv"
  `include "i2c_m_sequencer.sv"
  `include "i2c_m_agent.sv"


endpackage


