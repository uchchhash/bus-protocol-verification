`include "spi_defines2.sv"
`include "spi_clgen2.sv"
`include "spi_shift2.sv"
`include "spi_top2.sv"

