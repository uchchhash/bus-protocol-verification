//-------- SPI Base Sequence for SS line 0 ------------------//
class spi_base_sequence0 extends uvm_sequence#(spi_sequence_item);

    // Factory Registration
    `uvm_object_utils(spi_base_sequence0)


    // Constructor
    function new(string name = "spi_base_sequence0");
        super.new(name);
     //   `uvm_info(get_type_name(), "------ spi_base_sequence0 Constructed ------", UVM_HIGH)
    endfunction

    // ----- SPI Signals ----- //
    bit [6:0] char_len;
    bit [2:0] mode;
    bit ie;

    task body();
        `uvm_info(get_type_name(), "------ spi_base_sequence0 Body Task Started  ------", UVM_MEDIUM)
        `uvm_info(get_type_name(), "------ spi_base_sequence0 Body Task Finished ------", UVM_MEDIUM)
    endtask

endclass


//-------- SPI Base Sequence for SS line 1 ------------------//
class spi_base_sequence1 extends uvm_sequence#(spi_sequence_item);

    // Factory Registration
    `uvm_object_utils(spi_base_sequence1)


    // Constructor
    function new(string name = "spi_base_sequence1");
        super.new(name);
     //   `uvm_info(get_type_name(), "------ spi_base_sequence1 Constructed ------", UVM_HIGH)
    endfunction

    // ----- SPI Signals ----- //
    bit [6:0] char_len;
    bit [1:0] mode;
    bit ie;
    
    task body();
        `uvm_info(get_type_name(), "------ spi_base_sequence1 Body Task Started  ------", UVM_MEDIUM)
        `uvm_info(get_type_name(), "------ spi_base_sequence1 Body Task Finished ------", UVM_MEDIUM)
    endtask

endclass

//-------- SPI Base Sequence for SS line 2 ------------------//
class spi_base_sequence2 extends uvm_sequence#(spi_sequence_item);

    // Factory Registration
    `uvm_object_utils(spi_base_sequence2)


    // Constructor
    function new(string name = "spi_base_sequence2");
        super.new(name);
     //   `uvm_info(get_type_name(), "------ spi_base_sequence2 Constructed ------", UVM_HIGH)
    endfunction

    // ----- SPI Signals ----- //
    bit [6:0] char_len;
    bit [1:0] mode;
    bit ie;
    
    task body();
        `uvm_info(get_type_name(), "------ spi_base_sequence2 Body Task Started  ------", UVM_MEDIUM)
        `uvm_info(get_type_name(), "------ spi_base_sequence2 Body Task Finished ------", UVM_MEDIUM)
    endtask

endclass


//-------- SPI Base Sequence for SS line 3 ------------------//
class spi_base_sequence3 extends uvm_sequence#(spi_sequence_item);

    // Factory Registration
    `uvm_object_utils(spi_base_sequence3)


    // Constructor
    function new(string name = "spi_base_sequence3");
        super.new(name);
     //   `uvm_info(get_type_name(), "------ spi_base_sequence3 Constructed ------", UVM_HIGH)
    endfunction

    // ----- SPI Signals ----- //
    bit [6:0] char_len;
    bit [1:0] mode;
    bit ie;
    
    task body();
        `uvm_info(get_type_name(), "------ spi_base_sequence3 Body Task Started  ------", UVM_MEDIUM)
        `uvm_info(get_type_name(), "------ spi_base_sequence3 Body Task Finished ------", UVM_MEDIUM)
    endtask

endclass


//-------- SPI Base Sequence for SS line 4 ------------------//
class spi_base_sequence4 extends uvm_sequence#(spi_sequence_item);

    // Factory Registration
    `uvm_object_utils(spi_base_sequence4)


    // Constructor
    function new(string name = "spi_base_sequence4");
        super.new(name);
     //   `uvm_info(get_type_name(), "------ spi_base_sequence4 Constructed ------", UVM_HIGH)
    endfunction

    // ----- SPI Signals ----- //
    bit [6:0] char_len;
    bit [1:0] mode;
    bit ie;
    
    task body();
        `uvm_info(get_type_name(), "------ spi_base_sequence4 Body Task Started  ------", UVM_MEDIUM)
        `uvm_info(get_type_name(), "------ spi_base_sequence4 Body Task Finished ------", UVM_MEDIUM)
    endtask

endclass



//-------- SPI Base Sequence for SS line 5 ------------------//
class spi_base_sequence5 extends uvm_sequence#(spi_sequence_item);

    // Factory Registration
    `uvm_object_utils(spi_base_sequence5)


    // Constructor
    function new(string name = "spi_base_sequence5");
        super.new(name);
     //   `uvm_info(get_type_name(), "------ spi_base_sequence5 Constructed ------", UVM_HIGH)
    endfunction

    // ----- SPI Signals ----- //
    bit [6:0] char_len;
    bit [1:0] mode;
    bit ie;
    
    task body();
        `uvm_info(get_type_name(), "------ spi_base_sequence5 Body Task Started  ------", UVM_MEDIUM)
        `uvm_info(get_type_name(), "------ spi_base_sequence5 Body Task Finished ------", UVM_MEDIUM)
    endtask

endclass

//-------- SPI Base Sequence for SS line 6 ------------------//
class spi_base_sequence6 extends uvm_sequence#(spi_sequence_item);

    // Factory Registration
    `uvm_object_utils(spi_base_sequence6)


    // Constructor
    function new(string name = "spi_base_sequence6");
        super.new(name);
     //   `uvm_info(get_type_name(), "------ spi_base_sequence6 Constructed ------", UVM_HIGH)
    endfunction

    // ----- SPI Signals ----- //
    bit [6:0] char_len;
    bit [1:0] mode;
    bit ie;
    
    task body();
        `uvm_info(get_type_name(), "------ spi_base_sequence6 Body Task Started  ------", UVM_MEDIUM)
        `uvm_info(get_type_name(), "------ spi_base_sequence6 Body Task Finished ------", UVM_MEDIUM)
    endtask

endclass

//-------- SPI Base Sequence for SS line 7 ------------------//
class spi_base_sequence7 extends uvm_sequence#(spi_sequence_item);

    // Factory Registration
    `uvm_object_utils(spi_base_sequence7)


    // Constructor
    function new(string name = "spi_base_sequence7");
        super.new(name);
     //   `uvm_info(get_type_name(), "------ spi_base_sequence7 Constructed ------", UVM_HIGH)
    endfunction

    // ----- SPI Signals ----- //
    bit [6:0] char_len;
    bit [1:0] mode;
    bit ie;
    
    task body();
        `uvm_info(get_type_name(), "------ spi_base_sequence7 Body Task Started  ------", UVM_MEDIUM)
        `uvm_info(get_type_name(), "------ spi_base_sequence7 Body Task Finished ------", UVM_MEDIUM)
    endtask

endclass







