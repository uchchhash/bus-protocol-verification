package apb_spi_reg_seq_pkg;

    // Standard UVM import & include:
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    import env_pkg::*;
    import spi_reg_pkg::*;
    import apb_agnt_pkg::*;
    import spi_agnt_pkg::*;
    import intr_agnt_pkg::*;



    `include "apb_spi_reg_seq_base.sv"


endpackage
