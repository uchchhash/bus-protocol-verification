package apb_agnt_pkg;

    `include "uvm_macros.svh"
    import uvm_pkg::*;
    
    `include "apb_sequence_item.sv"
    `include "apb_base_sequence.sv"

    `include "apb_reset_sequence.sv"
    `include "apb_write_sequence.sv"
    `include "apb_read_sequence.sv"
   // `include "apb_random_sequence.sv"

    `include "apb_agent_config.sv"
    `include "apb_monitor.sv"
    `include "apb_driver.sv"
    `include "apb_sequencer.sv"
    `include "apb_agent.sv"
    `include "apb2reg_adapter.sv"


endpackage
