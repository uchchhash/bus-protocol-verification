package ahb_agnt_pkg;

	`include "uvm_macros.svh"
	 import uvm_pkg::*;


    `include "ahb_sequence_item.sv"
    `include "ahb_base_sequence.sv"
    `include "ahb_reset_sequence.sv"
    `include "ahb_write_sequence.sv"
    `include "ahb_read_sequence.sv"
    `include "ahb_random_sequence.sv"


    `include "ahb_sequencer.sv"
    `include "ahb_monitor.sv"
    `include "ahb_driver.sv"
    `include "ahb_coverage.sv"
    `include "ahb_agent_config.sv"
    `include "ahb_agent.sv"



endpackage
