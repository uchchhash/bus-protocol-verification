class testclass;


function testprint;
endfunct
