package env_pkg;

	`include "uvm_macros.svh"
	import uvm_pkg::*;
    import ahb_agnt_pkg::*;

    `include "ahb_predictor.sv"
    `include "scoreboard.sv"
    `include "environment_config.sv"
    `include "environment.sv"



endpackage
