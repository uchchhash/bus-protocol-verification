package agent_package;

	`include "uvm_macros.svh"
	import uvm_pkg::*;

	`include "ahb_sequence_item.sv"
	`include "ahb_sequence.sv"
	`include "ahb_sequencer.sv"
	`include "monitor.sv"
	`include "driver.sv"
	`include "ahb_coverage.sv"
	`include "agent_config.sv"
	`include "agent.sv"

endpackage
