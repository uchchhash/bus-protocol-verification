package apb_spi_test_seq_pkg;

    // Standard UVM import & include:
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    // Any further package imports:
    import apb_spi_reg_seq_pkg::*;
    import env_pkg::*;
    import spi_reg_pkg::*;
    import apb_agnt_pkg::*;
    import spi_agnt_pkg::*;
    import intr_agnt_pkg::*;



    // Includes:
    `include "apb_spi_vseq_base.sv"


endpackage
