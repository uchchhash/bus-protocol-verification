// This is a top level block.
// This block instantiates following blocks
// a) EgSlaveWIf
// b) EgSlaveRIf
// c) EgSlaveFn
// d) EgSlaveCIf

`include "EgSlaveAxi.v"

