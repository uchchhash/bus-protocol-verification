package environment_package;

	`include "uvm_macros.svh"
	import uvm_pkg::*;
	import agent_package::*;
	
	
    `include "scoreboard.sv"
    `include "environment_config.sv"
	`include "environment.sv"

endpackage
