
`include "timescale.v"
`include "timescale.v"
`include "i2cSlave_define.v"
`include "serialInterface.v"
`include "registerInterface.v"
`include "i2cSlave.v"
`include "i2cSlaveTop.v"
