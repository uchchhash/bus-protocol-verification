package agent_package;

	`include "uvm_macros.svh"
	 import uvm_pkg::*;

//	`include "apb_sequence_item.sv"
//	`include "apb_sequence.sv"
//	`include "apb_sequencer.sv"
//	`include "apb_monitor.sv"
//	`include "apb_driver.sv"
//	`include "coverage.sv"
//	`include "agent_config.sv"
//	`include "agent.sv"

endpackage
